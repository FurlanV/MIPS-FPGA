library verilog;
use verilog.vl_types.all;
entity divisorFrequencia is
    port(
        clk             : in     vl_logic;
        clock           : out    vl_logic
    );
end divisorFrequencia;
