module BANCOREGS(
input wire[4:0] rRegister1,
input wire[4:0] rRegister2,
input wire[4:0] writeRegister,
input wire[31:0] data,
input wire EscreveReg,
output wire[31:0] DadosLeitura1,
output wire[31:0] DadosLeitura2
);

 reg[31:0] registers[0:31];
 reg[31:0] temp1;
 reg[31:0] temp2;
 reg[31:0] tempWrite;
 
 
 initial
 begin
 
 registers[0] = 32'b00000000000000000000000000000000;
 registers[1] = 32'b00000000000000000000000000000000;
 registers[2] = 32'b00000000000000000000000000000000;
 registers[3] = 32'b00000000000000000000000000000000;
 registers[4] = 32'b00000000000000000000000000000000;
 registers[5] = 32'b00000000000000000000000000000000;
 registers[6] = 32'b00000000000000000000000000000000;
 registers[7] = 32'b00000000000000000000000000000000;
 registers[8] = 32'b00000000000000000000000000000101; //T0 = 5
 registers[9] = 32'b00000000000000000000000000000100; //T1 = 4
 registers[10] = 32'b0000000000000000000000000000101; //T2 = 5
 registers[11] = 32'b0000000000000000000000000000100; //T3 = 4
 registers[12] = 32'b00000000000000000000000000010000;
 registers[13] = 32'b00000000000000000000000001110000;
 registers[14] = 32'b00000000000000000000000011111111;
 registers[15] = 32'b00000000000000000000000000000111;
 registers[16] = 32'b00000000000000000000000000000010;
 registers[17] = 32'b00000000000000000000000000000001;
 registers[18] = 32'b00000000000000000000000000000001;
 registers[19] = 32'b00000000000000000000000000000000;
 registers[20] = 32'b00000000000000000000000000000000;
 registers[21] = 32'b00000000000000000000000000000000;
 registers[22] = 32'b00000000000000000000000000000000;
 registers[23] = 32'b00000000000000000000000000000000;
 registers[24] = 32'b00000000000000000000000000000000;
 registers[25] = 32'b00000000000000000000000000000000;
 registers[26] = 32'b00000000000000000000000000000000;
 registers[27] = 32'b00000000000000000000000000000000;
 registers[28] = 32'b00000000000000000000000000000000;
 registers[29] = 32'b00000000000000000000000000000000;
 registers[30] = 32'b00000000000000000000000000000000;
 registers[31] = 32'b00000000000000000000000000000000;
  
 end

 always @(rRegister1 or rRegister2)
 begin
 
 temp1 <= registers[rRegister1];
 temp2 <= registers[rRegister2];
 
 end

 always @(posedge EscreveReg)
 begin
 
 registers[writeRegister] <= data;
 
 end
 
 assign DadosLeitura1 = temp1;
 assign DadosLeitura2 = temp2;
 

endmodule